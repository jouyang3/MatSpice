This is a netlist		$must have a title line

r1	in	out	1000	$resistor connecting node 1 and 2
r2  out   3   500 $resistor
r3  out   0   250
v1  in   0   dc  6   $voltage source
.end				$Must have an end
